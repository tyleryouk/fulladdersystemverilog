module rc_adder_slice (
   // COMPLETE
);

    logic p, g;

    assign p = a ^ b;
    assign g = a & b;

    assign s     = // COMPLETE
    assign c_out = //COMPLETE

endmodule