module rc_adder4 (
 //COMPLETE
);

    logic [3:0] c;

    rc_adder_slice // COMPLETE USING ARRAY INSTANCING

    assign c[0] = // COMPLETE
    assign co = // COMPLETE

endmodule